/**
*
	*  des : regmaper
	*
	*
	*
*/

module macroreg #(

)(



);


endmodule 
