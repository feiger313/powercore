//==============================================
//   Filename       :
//   Author         :liuxf
//   Description    :
//   Called by      :
//   History        :
//   Email          :liuxf000@163.com
//   Company        :xxxx
//   Copyright(c) 2018,xxxx Technology Inc,All right reserved
//
//   //==============================================
//   

module fsm (



)


always @ (posedge mclk or negedge mreset_n)
begin
    if (!mreset_n)
	    test_reg   <= 1'b0 ;
    else
	    test_reg   <= 
end

endmodule
