//==============================================
//   Filename       :
//   Author         :liuxf
//   Description    :
//   Called by      :
//   History        :
//   Email          :liuxf000@163.com
//   Company        :xxxx
//   Copyright(c) 2018,xxxx Technology Inc,All right reserved
//
//   //==============================================
//   

module fsm (



)


endmodule
